// 用位掩码实现多路选择器
module mux5_8b (  
    input  [7:0]  in0, in1, in2, in3 ,in4,
    input  [2:0]  sel,
    output [7:0]  out 
);
assign out = ({8{sel==3'd0}} & in0)
           | ({8{sel==3'd1}} & in1)
           | ({8{sel==3'd2}} & in2)
           | ({8{sel==3'd3}} & in3)
           | ({8{sel==3'd4}} & in4)
endmodule
/*
这段代码使用了条件表达式和位掩码来实现多路选择器。我们逐部分分析：

{8{sel==3'd0}}：这是一个重复的位选择表达式，它会根据 sel==3'd0 的结果生成一个 8 位的掩码。如果 sel 等于 0，这个表达式的结果将是 8'b11111111（全 1）；否则，结果为 8'b00000000（全 0）。
& in0：将上面生成的 8 位掩码与 in0 进行按位与运算。只有当 sel 为 0 时，这个操作才会把 in0 的值传递到 out。
其他输入信号 in1、in2、in3 和 in4 的处理方式与 in0 类似。只有当 sel 等于相应的值时，对应的输入信号才会通过按位与运算传递到输出 out。
4. 按位选择
最终，所有的条件语句通过按位或（|）操作结合在一起。每个选择条件只会影响 out 的一部分，确保 out 的值只来自一个输入信号。换句话说，out 只会接收到与 sel 匹配的输入信号的值，而其他输入会被 "屏蔽"。

5. 工作原理
当 sel == 3'd0 时，out 仅等于 in0。
当 sel == 3'd1 时，out 仅等于 in1，其他输入（in0, in2, in3, in4）被屏蔽。
同理，其他值的 sel 会选择相应的输入信号。
*/